// Hi team, 
// Mic check 1, 2, 3. 

// Github is working? 